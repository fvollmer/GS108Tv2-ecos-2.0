# ====================================================================
#
#      io_flash.cdl
#
#      eCos IO configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      gthomas
# Original data:  gthomas
# Contributors:
# Date:           2000-07-06
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_IO_FLASH {
    display       "FLASH device drivers"
    include_dir   cyg/io
    description   "
        This option enables drivers for basic I/O services on
        flash devices."
    requires CYGPKG_ISOINFRA
    requires CYGINT_ISO_STRING_STRFUNCS

    compile       flash.c
 
    define_proc {
        puts $::cdl_header "#include <pkgconf/system.h>"
        puts $::cdl_header "#ifdef CYGDAT_IO_FLASH_DEVICE_HEADER"
        puts $::cdl_header "# include CYGDAT_IO_FLASH_DEVICE_HEADER"
        puts $::cdl_header "#endif "
    }

    cdl_option CYGNUM_FLASH_WORKSPACE_SIZE {
        display       "Extra memory required by FLASH device drivers"
	flavor        data
        default_value 0x1000
        description   "
            Use this option to control how much extra memory is used
            by the FLASH drivers to perform certain operations. This
            memory is used to hold driver functions in RAM (for platforms
            which require it).  The value should thus be large enough
            to hold any such driver.  Reducing this value will make
            more RAM available to general programs."
    }

    cdl_interface CYGHWR_IO_FLASH_DEVICE {
        display       "Hardware FLASH device drivers"
        description   "
            This option enables the hardware device drivers
            for the current platform."
    }

    cdl_interface CYGHWR_IO_FLASH_DEVICE_NOT_IN_RAM {
        display       "Hardware FLASH device drivers are not in RAM"
        flavor        booldata
        description   "
            This option makes the IO driver copy the device
            driver functions to RAM before calling them. Newer
            drivers should make sure that the functions are
            linked to RAM by putting them in .2ram sections."
    }

    cdl_interface CYGHWR_IO_FLASH_BLOCK_LOCKING {
        display       "Hardware can support block locking"
        flavor        booldata
        description   "
            This option will be enabled by devices which can support
            locking (write-protection) of individual blocks."
    }

    cdl_option CYGSEM_IO_FLASH_VERIFY_PROGRAM {
        display          "Verify data programmed to flash"
        flavor           bool
        default_value    1
        description      "
           Selecting this option will cause verification of data
           programmed to flash."
    }
    cdl_option CYGSEM_IO_FLASH_SOFT_WRITE_PROTECT {
        display          "Platform has flash soft DIP switch write-protect"
        flavor           bool
        default_value    0
        description      "
           Selecting this option will cause the state of a hardware jumper or
           dipswitch to be read by software to determine whether the flash is
           write-protected or not."
    }
    cdl_component CYGPKG_IO_FLASH_BLOCK_DEVICE {
        display         "Instantiate in I/O block device API"
        flavor          bool
        active_if       CYGPKG_IO
        default_value   0
        compile         -library=libextras.a flashiodev.c
        description     "
                Provides a block device accessible using the standard I/O
                API ( cyg_io_read() etc. )"

        cdl_component CYGDAT_IO_FLASH_BLOCK_DEVICE_NAME_1 {
                display       "Name of flash device 1 block device"
                flavor        data
                default_value { "\"/dev/flash1\"" }

            cdl_option CYGNUM_IO_FLASH_BLOCK_OFFSET_1 {
                display         "Start offset from flash base"
                flavor          data
                default_value   0x80000 
                description     "
                    This gives the offset from the base of flash which this
                    block device corresponds to."
            }
            cdl_option CYGNUM_IO_FLASH_BLOCK_LENGTH_1 {
                display         "Length"
                flavor          data
                default_value   0x1A0000
                description     "
                    This gives the length of the region of flash given over
                    to this block device."
            }
            
        }
                cdl_component CYGDAT_IO_FLASH_BLOCK_DEVICE_NAME_2 {
                display       "Name of flash device 1 block device"
                flavor        data
                default_value { "\"/dev/flash2\"" }

            cdl_option CYGNUM_IO_FLASH_BLOCK_OFFSET_2 {
                display         "Start offset from flash base"
                flavor          data
                default_value   0x220000 
                description     "
                    This gives the offset from the base of flash which this
                    block device corresponds to."
            }
            cdl_option CYGNUM_IO_FLASH_BLOCK_LENGTH_2 {
                display         "Length"
                flavor          data
                default_value   0x1A0000
                description     "
                    This gives the length of the region of flash given over
                    to this block device."
            }

        }
            cdl_component CYGDAT_IO_FLASH_BLOCK_DEVICE_NAME_3 {
                display       "Name of flash device 1 block device"
                flavor        data
                default_value { "\"/dev/boot.dim\"" }

            cdl_option CYGNUM_IO_FLASH_BLOCK_OFFSET_3 {
                display         "Start offset from flash base"
                flavor          data
                default_value   0x74000 
                description     "
                    This gives the offset from the base of flash which this
                    block device corresponds to."
            }
            cdl_option CYGNUM_IO_FLASH_BLOCK_LENGTH_3 {
                display         "Length"
                flavor          data
                default_value   0x8000
                description     "
                    This gives the length of the region of flash given over
                    to this block device."
            }

        }
               cdl_component CYGDAT_IO_FLASH_BLOCK_DEVICE_NAME_4 {
                display       "Name of flash device 4 block device"
                flavor        data
                default_value { "\"/dev/cfe\"" }

            cdl_option CYGNUM_IO_FLASH_BLOCK_OFFSET_4 {
                display         "Start offset from flash base"
                flavor          data
                default_value   0x000 
                description     "
                    This gives the offset from the base of flash which this
                    block device corresponds to."
            }
            cdl_option CYGNUM_IO_FLASH_BLOCK_LENGTH_4 {
                display         "Length"
                flavor          data
                default_value   0x80000
                description     "
                    This gives the length of the region of flash given over
                    to this block device."
            }

        }


    }
}
