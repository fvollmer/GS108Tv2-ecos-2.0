# ====================================================================
#
#      hal_mips_bcm53000.cdl
#
#      MIPS/BCM53000 variant architectural HAL package configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      
# Original data:  
# Contributors:
# Date:           
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_MIPS_BCM53000_BE {
    display       "MIPS BCM53000 variant HAL"
    parent        CYGPKG_HAL_MIPS
    hardware
    include_dir   cyg/hal
    define_header hal_mips_bcm53000.h
    description   "
           The BCM53000 variant HAL package provides generic support
           for platforms based on this variant. It is also necessary to
           select a specific target platform HAL package."

        cdl_option CYGHWR_HAL_MIPS_FPU {
            display    "Variant FPU support"
            calculated 0
        }

	cdl_option CYGPKG_HAL_MIPS_MSBFIRST {
            display    "CPU Variant little-endian"
            calculated 1
        }


    implements    CYGINT_HAL_MIPS_VARIANT    

    define_proc {
        puts $::cdl_header "#include <pkgconf/hal_mips.h>"
    }

    cdl_option CYGHWR_HAL_MIPS_CPU_FREQ_ACTUAL {
        display       "Actual CPU frequency"
        flavor        data
        legal_values  200000000 400000000
        default_value 400000000
        description "
            Only the frequency 200MHz is supported for this
            CPU variant."
    } 


    compile       var_misc.c var_intr.c

    make {
        <PREFIX>/lib/target.ld: <PACKAGE>/src/mips_bcm53000_be.ld
        $(CC) -E -P -Wp,-MD,target.tmp -DEXTRAS=1 -xc $(INCLUDE_PATH) $(CFLAGS) -o $@ $<
        @echo $@ ": \\" > $(notdir $@).deps
        @tail +2 target.tmp >> $(notdir $@).deps
        @echo >> $(notdir $@).deps
        @rm target.tmp
    }

    cdl_option CYGBLD_LINKER_SCRIPT {
        display "Linker script"
        flavor data
	no_define
        calculated  { "src/mips_bcm53000_be.ld" }
    }

    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        parent  CYGPKG_NONE
        description   "
	    Global build options including control over
	    compiler flags, linker flags and choice of toolchain."


        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { "mipsisa32-elf" }
            description "
                This option specifies the command prefix used when
                invoking the build tools."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
            default_value { "-mips32 -Wpointer-arith -Wstrict-prototypes -Winline -Wundef -Woverloaded-virtual -EB -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -fvtable-gc -finit-priority -fno-builtin -G0" }
            description   "
                This option controls the global compiler flags which
                are used to compile all packages by
                default. Individual packages may define
                options which override these global flags."
        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            default_value { "-mips32 -EB -nostdlib -Wl,--gc-sections -Wl,-static" }
            description   "
                This option controls the global linker flags. Individual
                packages may define options which override these global flags."
        }
    }
}

# EOF hal_mips_idt32334.cdl
