# ====================================================================
#
#      flash_mips_bcm947xx.cdl
#
#      FLASH memory - Flash memory support for BCM947xx boards
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
## Copyright (C) 2002 Gary Thomas
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      
# Contributors:   
# Date:           
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_FLASH_MIPS_BCM947xx {
    display       "FLASH memory support for BCM947xx boards"

    parent        CYGPKG_IO_FLASH
    active_if	  CYGPKG_IO_FLASH
    requires	  { CYGPKG_HAL_MIPS_BCM947xx || CYGPKG_HAL_MIPS_BCM953710}

    implements    CYGHWR_IO_FLASH_DEVICE

    include_dir   cyg/io

    compile       

    cdl_interface  CYGINT_DEVS_FLASH_CFI_REQUIRED {
        display    "CFI Flash driver required"
    }

    implements     CYGINT_DEVS_FLASH_CFI_REQUIRED

    define_proc {
        puts $::cdl_system_header "#define CYGDAT_DEVS_FLASH_CFI_CFG <cyg/io/flash_bcm947xx.h>"
        puts $::cdl_system_header "#define CYGDAT_DEVS_FLASH_JAG_CFG <cyg/io/flashDrvLib.h>"
    }

    compile   bcm947xx_flash.c nvram.c nvram_ecos.c flashDrvLib.c flash28f320DrvLib.c flash29lxxxDrvLib.c flash29GLxxxDrvLib.c flash28fxxxP33DrvLib.c
}
