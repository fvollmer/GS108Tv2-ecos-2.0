# ====================================================================
#
#      mips_bcm953000_et_drivers.cdl
#
#      Ethernet drivers - support for broadcom BCM953000 ethernet
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):     
# Contributors:  
# Date:          
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_ETH_BCM953000_ET_BE {
    display       "BCM953000 ethernet driver"
    description   "Ethernet driver for AMD PCNET compatible controllers."

    parent        CYGPKG_IO_ETH_DRIVERS
    active_if	  CYGPKG_IO_ETH_DRIVERS
    active_if     CYGPKG_HAL_MIPS_BCM953000_BE

    include_dir   cyg/devs/eth
    compile       -library=libextras.a etc.c et_ecos.c etcgmac.c
    # etc_adm.c

    define_proc {
        puts $::cdl_header "#include <pkgconf/system.h>";
	puts $::cdl_system_header \
       "#define CYGBLD_DEVS_ET_DEVICE_H <pkgconf/devs_eth_bcm953000_et_be.h>"
    }

    cdl_component CYGPKG_DEVS_ETH_ET0 {
        display       "ethernet port 0 driver"
        flavor        bool
        default_value 1

        implements CYGHWR_NET_DRIVERS
        implements CYGHWR_NET_DRIVER_ETH0
    }
    
    cdl_component CYGPKG_DEVS_ETH_ET1 {
        display       "ethernet port 1 driver"
        flavor        bool
        default_value 1

        implements CYGHWR_NET_DRIVERS
        implements CYGHWR_NET_DRIVER_ETH1
    }	
    
    cdl_option CYGNUM_DEVS_ETH_ET_DEV_COUNT {
	display "Number of supported interfaces."
	calculated    { 2 }
        flavor        data
	description   "
	    This option selects the number of PCI ethernet interfaces to
            be supported by the driver."
    }

    cdl_component CYGPKG_DEVS_ETH_BCM953000_ET_OPTIONS {
        display "BCM953000 ethernet driver build options"
        flavor  none
	no_define

        cdl_option CYGPKG_DEVS_ETH_BCM953000_ET_BE_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D_KERNEL -D__ECOS -DBCM47XX_CHOPS -DBCMDRIVER -I$(PREFIX)/include/cyg/hal/proto" }
            description   "
                This option modifies the set of compiler flags for
                building the BCM953000 ethernet driver
                package. These flags are used in addition to the set of
                global flags."
        }
    }
}
